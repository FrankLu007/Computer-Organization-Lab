//Subject:      CO project 3 - Shift_Left_Two_32
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer: 0416024 ������ 0516310 �f�ӿ�
//--------------------------------------------------------------------------------
//Date:        2017/5/12 11:42
//--------------------------------------------------------------------------------
//Description: Shift a 26bit number to the left by 2 bits
//  Output 28bit number
//--------------------------------------------------------------------------------

module Shift_Left_Two_28(
    data_i,
    data_o
    );

//I/O ports
input [26-1:0] data_i;
output [28-1:0] data_o;

//shift left 2

assign data_o[27:2] = data_i[25:0];
assign data_o[1:0] = 0;
endmodule
